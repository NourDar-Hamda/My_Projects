*** SPICE deck for cell NorGate{lay} from library Project
*** Created on Mon May 29, 2023 22:25:46
*** Last revised on Mon May 29, 2023 22:43:54
*** Written on Mon May 29, 2023 22:44:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NorGate{lay}
Mnmos@0 OUT IN1 gnd gnd nMos L=0.4U W=2.4U AS=5.52P AD=2.32P PS=13.2U PD=5.133U
Mnmos@1 gnd IN2 OUT gnd nMos L=0.4U W=2.4U AS=2.32P AD=5.52P PS=5.133U PD=13.2U
Mpmos@0 net@3 IN1 vdd vdd pMos L=0.4U W=2.4U AS=7.92P AD=1.2P PS=19U PD=3.4U
Mpmos@1 OUT IN2 net@3 vdd pMos L=0.4U W=2.4U AS=1.2P AD=2.32P PS=3.4U PD=5.133U

* Spice Code nodes in cell cell 'NorGate{lay}'
vdd VDD 0 DC 1.1
vin IN1 0 PULSE(0 1.1 0n 1n 1n 20n 40n 10)
vin1 IN2 0 PULSE(0 1.1 0n 1n 1n 40n 80n 10)
cload OUT 0 5fF
.tran 0 160n
.include C:\Users\NOR0185869\Downloads\Tech_models.txt
.END
.END
