*** SPICE deck for cell InvGate{lay} from library Project
*** Created on Mon May 29, 2023 21:25:19
*** Last revised on Mon May 29, 2023 21:50:20
*** Written on Mon May 29, 2023 21:51:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: InvGate{lay}
Mnmos@0 OUT IN gnd gnd nMos L=0.4U W=2.4U AS=7.92P AD=3.12P PS=19U PD=7.4U
Mpmos@0 OUT IN vdd vdd pMos L=0.4U W=2.4U AS=7.32P AD=3.12P PS=17.8U PD=7.4U

* Spice Code nodes in cell cell 'InvGate{lay}'
vdd VDD 0 DC 1.1
vin IN 0 PULSE(0 1.1 0n 1n 1n 20n 40n 10)
cload OUT 0 0fF
.tran 0 160n
.include C:\Users\NOR0185869\Downloads\Tech_models.txt
.END
.END
